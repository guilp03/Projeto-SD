module timer_controle(keypad, enablen, clk100, D, loadn, pgt_1Hz);
        input wire [9:0] keypad;
        input wire enablen clk100;
        output wire [3:0] D;
        output wire loadn, pgt_1Hz;
endmodule