$date
	Mon Oct 17 12:41:09 2022
$end
$version
	Icarus Verilog
$end
$timescale
	1ns
$end
$scope module control_mag_teste $end
$var wire 1 ! reset_TB $end
$var wire 1 " set_TB $end
$var reg 1 # clearn_TB $end
$var reg 1 $ door_closed_TB $end
$var reg 1 % startn_TB $end
$var reg 1 & stopn_TB $end
$var reg 1 ' timer_done_TB $end
$scope module DUT $end
$var wire 1 ( clearn $end
$var wire 1 ) door_closed $end
$var wire 1 * startn $end
$var wire 1 + stopn $end
$var wire 1 , timer_done $end
$var reg 1 - reset $end
$var reg 1 . set $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
x.
1-
0,
0+
1*
0)
0(
0'
0&
1%
0$
0#
x"
1!
$end
#5
0-
0!
1.
1"
1$
1)
#10
1-
1!
1&
1+
#15
0-
0!
0&
0+
#20
1-
1!
1'
1,
#25
0'
0,
0$
0)
#30
1'
1,
1$
1)
1#
1(
#35
0-
0!
0'
0,
0#
0(
#40
1-
1!
1'
1,
1#
1(
1&
1+
#45
0%
0*
#50
0'
0,
0$
0)
0#
0(
0&
0+